// desgin constant

// topmodule
`define PERSON_COUNTER_DATA_WIDTH                   16

`define COMMAND_CONTROL_TYPE_WIDTH                  3
`define COMMAND_CONTROL_DATA_WIDTH                  8

`define HOME_WINDOW_COUNT                           8
`define HOME_DOOR_COUNT                             4

`define TEMPERATURE_SENSOR_DATA_WIDTH               8
`define TEMPERATURE_SENSOR_MIN_TEMP                 7 // 7 derece altına düşerse ISIT
`define TEMPERATURE_SENSOR_MAX_TEMP                 20 // 20 derece altına düşerse SOĞUT
`define AC_COOL_MODE_BIT                            0
`define AC_HEAT_MODE_BIT                            1
