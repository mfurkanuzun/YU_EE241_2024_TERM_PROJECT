// desgin constant

// topmodule
`define PERSON_COUNTER_DATA_WIDTH                   16


`define HOME_WINDOW_COUNT                           8
`define HOME_DOOR_COUNT                             4

`define TEMPERATURE_SENSOR_DATA_WIDTH               8

