`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.11.2024 20:10:02
// Design Name: 
// Module Name: security_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "design_constant.vh"

module security_controller
    (
        input [`PERSON_COUNTER_DATA_WIDTH-1:0] person_count_i
    );
endmodule



















